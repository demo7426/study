/*************************************************
Copyright (C), 2009-2012    , Level Chip Co., Ltd.
�ļ���:	tb_led.v
��  ��:	Ǯ��      �汾: V0.1.0     �½�����: 2025.11.27
��  ��: ʵ�ֶ�led��ˮ�ƵĲ���
��  ע:	
�޸ļ�¼:

  1.  ����: 2025.11.27
      ����: Ǯ��
      ����:
          1) ��Ϊģ���һ���汾��
      �汾:V0.1.0

*************************************************/

`timescale 1ns/1ns      //���浥λ/���澫��

module tb_flow_led();

parameter CLK_PERIOD = 20;  //ʱ������20ns

reg sys_clk;
reg sys_rst_n;

wire [1:0] led;

//�źų�ʼ��
initial begin
    sys_clk <= 1'b0;
    sys_rst_n <= 1'b0;
    #200
    sys_rst_n <= 1'b1;
end

//����ʱ��
always #(CLK_PERIOD/2) sys_clk = ~sys_clk;

//�����������
flow_led u_flow_led(
    .sys_clk        (sys_clk),
    .sys_rst_n      (sys_rst_n),
    .led            (led)
    );

endmodule