/*************************************************
Copyright (C), 2009-2012    , Level Chip Co., Ltd.
�ļ���:	led.v
��  ��:	Ǯ��      �汾: V0.1.0     �½�����: 2025.06.02
��  ��: ����led��
��  ע:	
�޸ļ�¼:

  1.  ����: 2025.06.02
      ����: Ǯ��
      ����:
          1) ��Ϊģ���һ���汾��
      �汾:V0.1.0

*************************************************/

module led (
    input key,      //���밴��,Ĭ��Ϊ�ߵ�ƽ
    output led      //���LED,�ߵ�ƽ����
);

//��key = 1, led = 0; ��key = 0, led = 1; 
assign led = ~key;
    
endmodule


