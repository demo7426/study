/*************************************************
Copyright (C), 2009-2012    , Level Chip Co., Ltd.
�ļ���:	tb_led.v
��  ��:	Ǯ��      �汾: V0.1.0     �½�����: 2025.06.02
��  ��: ʵ�ֶԵ���led�ƵĲ���
��  ע:	
�޸ļ�¼:

  1.  ����: 2025.06.02
      ����: Ǯ��
      ����:
          1) ��Ϊģ���һ���汾��
      �汾:V0.1.0

*************************************************/

`timescale 1ns/1ns      //��λ/����

module tb_led();

reg key;
wire led;

initial begin
     key <= 1'b1;
     #200
     key <= 1'b0;
     #500
     key <= 1'b1;
     #1000
     key <= 1'b0;
     #1000
     key <= 1'b1;    
end

led u_led(
    .key (key),
    .led (led)
);

endmodule